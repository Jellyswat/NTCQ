** Profile: "SCHEMATIC1-123"  [ e:\����\2018-2019ũ���������Ŀ\��ѹ&di_dv\didv-pspicefiles\schematic1\123.sim ] 

** Creating circuit file "123.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "d:/ddd/213/opa4330_pspice_aio/opa4330.lib" 
* From [PSPICE NETLIST] section of E:\BaiduNetdisk\Cadence\Cadence\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 5u 0 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END

** Profile: "SCHEMATIC1-ex1"  [ C:\Users\wxy\Desktop\��Ŀ����\��Ŀ����\��ֵ���ֵ�·�������\��Ŀ2016(��ֵ��\pspice\ex1\ex1-pspicefiles\schematic1\ex1.sim ] 

** Creating circuit file "ex1.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of F:\8848\Cadence\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 1 0 1m 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END

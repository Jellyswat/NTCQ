** Profile: "SCHEMATIC1-nwe"  [ D:\ddd\gkd\2018-2019ũ���������Ŀ\RCC���ص�Դ2.0\111-pspicefiles\schematic1\nwe.sim ] 

** Creating circuit file "nwe.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of F:\8848\Cadence\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 500m 0 SKIPBP 
.OPTIONS ADVCONV
.OPTIONS ABSTOL= 1p
.OPTIONS GMIN= 1p
.OPTIONS VNTOL= 1u
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END

** Profile: "SCHEMATIC1-nwe"  [ G:\BaiduNetdiskDownload\����\2018-2019ũ���������Ŀ\RCC���ص�Դ1.0\111-pspicefiles\schematic1\nwe.sim ] 

** Creating circuit file "nwe.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of E:\BaiduNetdisk\Cadence\Cadence\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 200u 0 SKIPBP 
.OPTIONS ADVCONV
.OPTIONS ABSTOL= 1p
.OPTIONS GMIN= 1p
.OPTIONS VNTOL= 1u
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END

** Profile: "SCHEMATIC1-6666"  [ D:\ddd\gkd\2018-2019ũ���������Ŀ\΢С����ת��pdf��·ͼ\heiheihei-pspicefiles\schematic1\6666.sim ] 

** Creating circuit file "6666.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of F:\8848\Cadence\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "E:\Cadence\SPB_17.2\tools\pspice\library\nom.lib" 

*Analysis directives: 
.DC LIN I_I1 0A 100nA 10nA 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
